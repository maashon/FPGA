`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
module DEC3to8();


endmodule
