`timescale 1ns / 1ps
module bus(sel,in,out);
input [2:0] sel;
input [15:0] in;
output [15:0] out;

//MEMORY mm();
//REGISTER12 AR(
//REGISTER12 PC(
//REGISTER DR(
//REGISTER IR(
//REGISTER TR(
//REGISTER AC(

endmodule
